// $Id: $
// File name:   sample.sv
// Created:     2/23/2021
// Author:      Rushabh Ranka
// Lab Section: 337-07
// Version:     1.0  Initial Design Entry
// Description: sample.
